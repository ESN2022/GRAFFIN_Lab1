
module Lab1_qsys (
	clk_clk,
	pio_0_export,
	rst_reset_n,
	pio_1_export);	

	input		clk_clk;
	output	[7:0]	pio_0_export;
	input		rst_reset_n;
	input		pio_1_export;
endmodule
